`ifndef __proc_defs
`define __proc_defs

`define NUM_THREADS 8

`endif
