

module rnd_mtcpu_tb();


endmodule